/*
   Arquitetura de Computadores I - Guia_04,

   Nome: Larissa Valadares Silqueira
   Matricula: 754065-5
*/

// expressao
module fxyz (output s1, s2, input x, y);
   assign s1 = ~(~y | x) & (~y | x);
   assign s2 = (y & ~x) & (~y | x);
endmodule

// teste
module test_module;

   reg x, y;
   wire se, ss;

   // instancias
   fxyz FXYZ (se, ss, x, y);

   // valores iniciais
   initial begin: start
      
      x = 1'b0;
      y = 1'b0;

   end

   // parte principal
   initial begin: main
      $display("-------- Guia0402-e --------\n");
   
      $display("e) (y' + x)' . (y' + x) = s\n   (y . x') . (y' + x) = ss\n\n   x y   s ss");
      $monitor("   %b %b = %b %b", x, y, se, ss);
      #1 x=0; y=0;
      #1 x=0; y=1;
      #1 x=1; y=0;
      #1 x=1; y=1;

   end

endmodule

/*

   -------- Guia0402-e --------

   e) (y' + x)' . (y' + x) = s
      (y . x') . (y' + x) = ss

      x y   s ss
      0 0 = 0 0
      0 1 = 0 0
      1 0 = 0 0
      1 1 = 0 0

*/
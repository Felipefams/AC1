// -------------------------
// Exemplo_0501 - GATES
// Nome: xxx yyy zzz
// Matricula: 999999
// -------------------------

// -------------------------
// f5_gate
// m a b s
// 0 0 0 0
// 1 0 1 1 <- a'.b
// 2 1 0 1 <- a ^ b
// 3 1 1 0
//
// -------------------------

module f5a ( output s,
    input a,
    input b );

    // definir dado local

    wire nor_a;
    wire nor_b;
    wire nor_c;
    wire nor_c2;
    

    // descrever por portas

    nor NOR1 ( nor_a, a, a );
    nor NOR2 ( nor_b, b, b );
    nor NOR3 ( nor_c, nor_a, nor_b );
    nor NOR4 ( nor_c2, a, b );
    nor NOR5 ( s, nor_c, nor_c2 );
    //and AND1 ( s, not_a, b );
endmodule // f5a

// -------------------------
// f5_gate
// m a b s
// 0 0 0 0
// 1 0 1 1 <- a ^ b
// 2 1 0 1 <- a ^ b
// 3 1 1 0
//
// -------------------------

module f5b ( output s,
input a,
input b );

// descrever por expressao

assign s = a ^ b;
endmodule // f5b

module test_f5;

    // ------------------------- definir dados

    reg x;
    reg y;
    wire a, b;
    f5a moduloA ( a, x, y );
    f5b moduloB ( b, x, y );

    // ------------------------- parte principal

    initial
    begin : main
        $display("Exemplo_0507 - MARCUS PRADO SILVA - 753117");
        $display("Test module");
        $display("   x     y     a     b");
        
        // projetar testes do modulo

        $monitor("%4b  %4b  %4b  %4b", x, y, a, b);
        x = 1'b0; y = 1'b0;
        #1 x = 1'b0; y = 1'b1;
        #1 x = 1'b1; y = 1'b0;
        #1 x = 1'b1; y = 1'b1;
    end
endmodule // test_f5
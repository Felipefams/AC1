// -------------------------
// Exemplo_0804 - 
// Nome:Felipe Augusto Morais Silva 
// Matricula:748473 
// -------------------------
// -------------------------
// 1's complement 
// -------------------------
module comp1 (output s, input a);
not NOT1(s, a);
endmodule // inequality operator
//full adder
module fullAdder ( output sum, output cout, input a, input b, input cin );
	assign {sum,cout} = a + b + cin;
endmodule // fullAdder
//2's complement
module comp2 (output sum, output cout, input a, input b, input carry);
	wire comp_1,comp_2;
	comp1(comp_1, a);
	comp1(comp_2, b);
	fullAdder(sum,cout, comp1, comp2, 1);
endmodule
module halfSubTeste;
reg a, b, carry;
carry = 1;
wire cout,sum;
comp2 teste(sum, cout, a, b, carry);
initial begin
$display("Exemplo0804 - Felipe Augusto Morais Silva- 748473");
$display("Test ALU's comp2 test");
$display("   a       b =   sum     cout");
$monitor("%6b    %6b = %6b    %6b", a, b, sum, cout);
           a = 6'b000000; b = 6'b000001; 
		#1 a = 6'b000000; b = 6'b000010; 
		#1 a = 6'b000000; b = 6'b000011; 
		#1 a = 6'b000000; b = 6'b000100; 
		#1 a = 6'b000000; b = 6'b000101; 
		#1 a = 6'b000000; b = 6'b000110; 
		#1 a = 6'b000000; b = 6'b000111; 
		#1 a = 6'b000000; b = 6'b010001; 
		#1 a = 6'b000000; b = 6'b010010; 
		#1 a = 6'b000000; b = 6'b010011; 
		#1 a = 6'b000000; b = 6'b010100; 
		#1 a = 6'b000000; b = 6'b101101; 
		#1 a = 6'b000000; b = 6'b101110; 
		#1 a = 6'b000000; b = 6'b101111; 
		#1 a = 6'b000000; b = 6'b110000; 
		#1 a = 6'b000000; b = 6'b110001; 
		#1 a = 6'b000000; b = 6'b110110; 
		#1 a = 6'b000000; b = 6'b110111; 
		#1 a = 6'b000000; b = 6'b111000; 
		#1 a = 6'b000000; b = 6'b111001; 
		#1 a = 6'b000000; b = 6'b111010; 
		#1 a = 6'b000000; b = 6'b111011; 
		#1 a = 6'b000000; b = 6'b111100; 
		#1 a = 6'b000000; b = 6'b111101; 
		#1 a = 6'b000000; b = 6'b111110; 
		#1 a = 6'b000000; b = 6'b111111; 

		#1 a = 6'b000010; b = 6'b111111; 
		#1 a = 6'b000011; b = 6'b111111; 
		#1 a = 6'b000100; b = 6'b111111; 
		#1 a = 6'b000101; b = 6'b111111; 
		#1 a = 6'b000110; b = 6'b111111; 
		#1 a = 6'b000111; b = 6'b111111; 
		#1 a = 6'b001000; b = 6'b111111; 
		#1 a = 6'b001001; b = 6'b111111; 
		#1 a = 6'b001010; b = 6'b111111; 
		#1 a = 6'b001011; b = 6'b111111; 
		#1 a = 6'b001100; b = 6'b111111; 
		#1 a = 6'b001101; b = 6'b111111; 
		#1 a = 6'b001110; b = 6'b111111; 
		#1 a = 6'b001111; b = 6'b111111; 
		#1 a = 6'b010000; b = 6'b111111; 
		#1 a = 6'b010001; b = 6'b111111; 
		#1 a = 6'b010010; b = 6'b111111; 
		#1 a = 6'b010011; b = 6'b111111; 
		#1 a = 6'b010100; b = 6'b111111; 
		#1 a = 6'b010101; b = 6'b111111; 
		#1 a = 6'b010110; b = 6'b111111; 
		#1 a = 6'b010111; b = 6'b111111; 
		#1 a = 6'b011000; b = 6'b111111; 
		#1 a = 6'b011001; b = 6'b111111; 
		#1 a = 6'b011010; b = 6'b111111; 
		#1 a = 6'b011011; b = 6'b111111; 
		#1 a = 6'b011100; b = 6'b111111; 
		#1 a = 6'b011101; b = 6'b111111; 
		#1 a = 6'b011110; b = 6'b111111; 
		#1 a = 6'b011111; b = 6'b111111; 
		#1 a = 6'b100000; b = 6'b111111; 
		#1 a = 6'b100001; b = 6'b111111; 
		#1 a = 6'b100010; b = 6'b111111; 
		#1 a = 6'b100011; b = 6'b111111; 
		#1 a = 6'b100100; b = 6'b111111; 
		#1 a = 6'b100101; b = 6'b111111; 
		#1 a = 6'b100110; b = 6'b111111; 
		#1 a = 6'b100111; b = 6'b111111; 
		#1 a = 6'b101000; b = 6'b111111; 
		#1 a = 6'b101001; b = 6'b111111; 
		#1 a = 6'b101010; b = 6'b111111; 
		#1 a = 6'b101011; b = 6'b111111; 
		#1 a = 6'b111110; b = 6'b111111; 
		#1 a = 6'b111111; b = 6'b111111; 

		#1 a = 6'b100010; b = 6'b100010; 
		#1 a = 6'b100011; b = 6'b100011; 
		#1 a = 6'b100100; b = 6'b100100; 
		#1 a = 6'b100101; b = 6'b100101; 
		#1 a = 6'b000001; b = 6'b000001; 
		#1 a = 6'b111111; b = 6'b111111; 
		#1 a = 6'b100010; b = 6'b100010; 
		#1 a = 6'b100011; b = 6'b100011; 
		#1 a = 6'b100100; b = 6'b100100; 
		#1 a = 6'b100101; b = 6'b100101; 
		#1 a = 6'b000001; b = 6'b000001; 
		#1 a = 6'b111111; b = 6'b111111; 

end
endmodule // test_fullAdder
